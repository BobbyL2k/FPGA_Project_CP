module uart_recevier(
  
);

endmodule // uart_recevier